//module p2interface(
//	input [9:0]  p2_PosX, p2_PosY, p2_SizeX, p2_SizeY,
//	input logic p2_in_air, p2_crouch, p2_move_right, p2_move_left, p2_dir, p2_kick, p2_punch,
//	input [2:0] p2_run_state
//);